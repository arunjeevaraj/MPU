-- normalize the input between 1<= x < 2 
-- Normalize value maps to a lookup table

library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

entity normal is
    port( clk : in std_logic;
	      rst : in std_logic;
	      data_diag : in std_logic_vector(31 downto 0);   --Diagonal elements as input
		  
		  o_norm : out std_logic_vector(10 downto 0); --Normalize value 
		  norm_sig : out std_logic_vector(1 downto 0);  --norm_sig is to determine how many bits required in de-normalization
	      o_xi : out std_logic_vector(15 downto 0)    -- Initial estimate based on normalize data
		  );
end normal;

architecture behav of normal is
signal temp : std_logic_vector(15 downto 0) := (others => '0');
signal temp_o_norm,i_div : std_logic_vector(10 downto 0) := (others => '0');
signal norm : std_logic := '0';

begin
i_div <= data_diag(18 downto 8);   --Taking 7 bits for fraction and 3 bits for interger,Total 10 bits
o_norm <= temp_o_norm;
process(clk)
begin
     if  rising_edge(clk) then
	    if rst = '1' then
		   temp_o_norm <= (others => '0');
		   norm <='0';
		   norm_sig <= "00";
	    elsif i_div(10)='1' and i_div(9)='1' then    --Normalize incoming data 1<= x<2 by shifting bits to right and set a flag for it
		   temp_o_norm <= "00" & i_div(10 downto 2);
		   norm <='1';
		   norm_sig <= "10";
		elsif i_div(10)='1' and i_div(9)='0' then 
		   temp_o_norm <= "00" & i_div(10 downto 2);
		   norm <='1';
		   norm_sig <= "10";
		elsif i_div(9) ='1' then
		   temp_o_norm <= '0' & i_div(10 downto 1);
		   norm <='1';
		   norm_sig <= "01";
		elsif data_diag(31)='1' then 
		   temp_o_norm <= i_div;
		   norm <= '1';
		   norm_sig <= "11";   --For sign bit
		else 
		   temp_o_norm <= i_div;
		   norm <= '1';
		   norm_sig <= "00";
		end if;
	end if;
end process;

lut : process(norm,temp_o_norm,temp)
begin
if norm='1' then
   o_xi <= temp;
   
else 
   o_xi <= (others => '0');
end if;
--LUT with 128 entries 
case temp_o_norm is 
    when "00010000000" =>
	      temp <= "1111000011100011";  
    when "00010000001" =>
	      temp <= "1111000011000110";   
	when "00010000010" =>
	      temp <= "1111000010101010";   
	when "00010000011" =>
	      temp <= "1111000010001110";   
	when "00010000100" =>
	      temp <= "1111000001110010";   
	when "00010000101" =>
	      temp <= "1111000001010101";   
	when "00010000110" =>
	      temp <= "1111000000111001";   
	when "00010000111" =>
	      temp <= "1111000000011101";   
	when "00010001000" =>
	      temp <= "1111000000000001";   
 	when "00010001001" =>
	      temp <= "1110111111100101";   
	when "00010001010" =>
	      temp <= "1110111111001001";   
	when "00010001011" =>
	      temp <= "1110111110101101";   
	when "00010001100" =>
	      temp <= "1110111110010001";   
	when "00010001101" =>
	      temp <= "1110111101110101";   
    when "00010001110" =>
	      temp <= "1110111101011001";   
    when "00010001111" =>
	      temp <= "1110111100111101";	   
    when "00010010000" =>
	      temp <= "1110111100100001";  
    when "00010010001" =>
	      temp <= "1110111100000101";   
	when "00010010010" =>
	      temp <= "1110111011101001";   
	when "00010010011" =>
	      temp <= "1110111011001101";   
	when "00010010100" =>
	      temp <= "1110111010110001";   
	when "00010010101" =>
	      temp <= "1110111010010101";   
	when "00010010110" =>
	      temp <= "1110111001111010";   
	when "00010010111" =>
	      temp <= "1110111001011110";   
	when "00010011000" =>
	      temp <= "1110111001000010";   
 	when "00010011001" =>
	      temp <= "1110111000100110";   
	when "00010011010" =>
	      temp <= "1110111000001011";   
	when "00010011011" =>
	      temp <= "1110110111101111";   
	when "00010011100" =>
	      temp <= "1110110111010100";   
	when "00010011101" =>
	      temp <= "1110110110111000";   
    when "00010011110" =>
	      temp <= "1110110110011100";   
    when "00010011111" =>
	      temp <= "1110110110000001";	   
    when "00010100000" =>
	      temp <= "1110110101100101";  
    when "00010100001" =>
	      temp <= "1110110101001010";   
	when "00010100010" =>
	      temp <= "1110110100101110";   
	when "00010100011" =>
	      temp <= "1110110100010011";   
	when "00010100100" =>
	      temp <= "1110110011110111";   
	when "00010100101" =>
	      temp <= "1110110011011100";   
	when "00010100110" =>
	      temp <= "1110110011000001";   
	when "00010100111" =>
	      temp <= "1110110010100101";   
	when "00010101000" =>
	      temp <= "1110110010001010";   
 	when "00010101001" =>
	      temp <= "1110110001101111";   
	when "00010101010" =>
	      temp <= "1110110001010011";   
	when "00010101011" =>
	      temp <= "1110110000111000";   
	when "00010101100" =>
	      temp <= "1110110000011101";   
	when "00010101101" =>
	      temp <= "1110110000000010";   
    when "00010101110" =>
	      temp <= "1110101111100110";   
    when "00010101111" =>
	      temp <= "1110101111001011";	   
    when "00010110000" =>
	      temp <= "1110101110110000";  
    when "00010110001" =>
	      temp <= "1110101110010101";   
	when "00010110010" =>
	      temp <= "1110101101111010";   
	when "00010110011" =>
	      temp <= "1110101101011111";   
	when "00010110100" =>
	      temp <= "1110101101000100";   
	when "00010110101" =>
	      temp <= "1110101100101001";   
	when "00010110110" =>
	      temp <= "1110101100001110";   
	when "00010110111" =>
	      temp <= "1110101011110011";   
	when "00010111000" =>
	      temp <= "1110101011011000";   
 	when "00010111001" =>
	      temp <= "1110101010111101";   
	when "00010111010" =>
	      temp <= "1110101010100010";   
	when "00010111011" =>
	      temp <= "1110101010000111";   
	when "00010111100" =>
	      temp <= "1110101001101100";   
	when "00010111101" =>
	      temp <= "1110101001010010";   
    when "00010111110" =>
	      temp <= "1110101000110111";   
    when "00010111111" =>
	      temp <= "1110101000011100";	   
    when "00011000000" =>
	      temp <= "1110101000000001";  
    when "00011000001" =>
	      temp <= "1110100111100111";   
	when "00011000010" =>
	      temp <= "1110100111001100";   
	when "00011000011" =>
	      temp <= "1110100110110001";   
	when "00011000100" =>
	      temp <= "1110100110010110";   
	when "00011000101" =>
	      temp <= "1110100101111100";   
	when "00011000110" =>
	      temp <= "1110100101100001";   
	when "00011000111" =>
	      temp <= "1110100101000111";   
	when "00011001000" =>
	      temp <= "1110100100101100";   
 	when "00011001001" =>
	      temp <= "1110100100010010";   
	when "00011001010" =>
	      temp <= "1110100011110111";   
	when "00011001011" =>
	      temp <= "1110100011011101";   
	when "00011001100" =>
	      temp <= "1110100011000010";   
	when "00011001101" =>
	      temp <= "1110100010101000";   
    when "00011001110" =>
	      temp <= "1110100010001101";   
    when "00011001111" =>
	      temp <= "1110100001110011";	   	
    when "00011010000" =>
	      temp <= "1110100001011000";   
	when "00011010001" =>
	      temp <= "1110100000111110";   
	when "00011010010" =>
	      temp <= "1110100000100100";   
	when "00011010011" =>
	      temp <= "1110100000001010";   
	when "00011010100" =>
	      temp <= "1110011111101111";   
	when "00011010101" =>
	      temp <= "1110011111010101";   
	when "00011010110" =>
	      temp <= "1110011110111011";   
 	when "00011010111" =>
	      temp <= "1110011110100001";   
	when "00011011000" =>
	      temp <= "1110011110000110";   
	when "00011011001" =>
	      temp <= "1110011101101100";   
	when "00011011010" =>
	      temp <= "1110011101010010";   
	when "00011011011" =>
	      temp <= "1110011100111000";   
    when "00011011100" =>
	      temp <= "1110011100011110";   
    when "00011011101" =>
	      temp <= "1110011100000100";	   	
    when "00011011110" =>
	      temp <= "1110011011101010";   
	when "00011011111" =>
	      temp <= "1110011011010000";   
	when "00011100000" =>
	      temp <= "1110011010110110";   
	when "00011100001" =>
	      temp <= "1110011010011100";   
	when "00011100010" =>
	      temp <= "1110011010000010";   
	when "00011100011" =>
	      temp <= "1110011001101000";   
	when "00011100100" =>
	      temp <= "1110011001001110";   
 	when "00011100101" =>
	      temp <= "1110011000110100";   
	when "00011100110" =>
	      temp <= "1110011000011010";   
	when "00011100111" =>
	      temp <= "1110011000000000";   
	when "00011101000" =>
	      temp <= "1110010111100111";   
	when "00011101001" =>
	      temp <= "1110010111001101";   
    when "00011101010" =>
	      temp <= "1110010110110011";   
    when "00011101011" =>
	      temp <= "1110010110011001";	   	
    when "00011101100" =>
	      temp <= "1110010101111111";   
	when "00011101101" =>
	      temp <= "1110010101100110";   
	when "00011101110" =>
	      temp <= "1110010101001100";   
	when "00011101111" =>
	      temp <= "1110010100110010";   
	when "00011110000" =>
	      temp <= "1110010100011001";   
	when "00011110001" =>
	      temp <= "1110010011111111";   
	when "00011110010" =>
	      temp <= "1110010011100110";   
 	when "00011110011" =>
	      temp <= "1110010011001100";   
	when "00011110100" =>
	      temp <= "1110010010110010";   
	when "00011110101" =>
	      temp <= "1110010010011001";   
	when "00011110110" =>
	      temp <= "1110010001111111";   
	when "00011110111" =>
	      temp <= "1110010001100110";   
    when "00011111000" =>
	      temp <= "1110010001001100";   
    when "00011111001" =>
	      temp <= "1110010000110011";	   	
    when "00011111010" =>
	      temp <= "1110010000011010";   
	when "00011111011" =>
	      temp <= "1110010000000000";   
	when "00011111100" =>
	      temp <= "1110001111100111";   
	when "00011111101" =>
	      temp <= "1110001111001110";   
	when "00011111110" =>
	      temp <= "1110001110110100";   
	when "00011111111" =>
	      temp <= "1110001110011011";   		  
	when others =>
	      temp <= "1110001110000010";
		  
end case;
end process;
end behav;


