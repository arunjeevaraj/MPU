-- File   : mat_ctrl.vhd
-- Author : Arun jeevaraj
-- Team   : Arun and Deepak Yadav  Team Mentor : Liang Liu 
-- usage  : level 2 of control flow , interfaces the address decoder and master controller. , has statemachines for all the modes of instructions
--			supported by master controller. generates the required control signals for data flow and address decoder.
-- DLM    : 6/23/2016   7:36 AM 
-- Tested : modelsim student edition 10.4 a
-- Todo   : removes ram_sel_stored with rs_ram_sel , it is redundant. 
-- error  : none.
-- warning: none. 
-- copyright : Arun Jeevaraj .c 2016 Lund University.

library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

---- A map of instruction to mode control signals that mat controller supports. 
-- mode 000 for loading the input matrix to ram, to op_r -- done
-- mode 001 for performing mat_mult. op_1*op_2 = op_r    -- doing now.
-- mode 010 for diag multiply operation spec_command = 000 --> diag to matrix  and spec_command= 001  --> matrix to diag mulitplication.
-- mode 011 for adding or subtraction identity matrix.     special command 000 for adding and special command 001 for subtraction.
-- mode 100 for mat copy --  op_1 to op_r.     
-- mode 101 -- reserved for matrix matrix addition.
-- mode 110 -- reserved for matrit matrix dot product.
-- mode 111 for sending the result out serially through data out col wise..


entity mat_ctrl_v1 is
port (
			start     : in std_logic; 								-- handshake signals
			done      : out std_logic;
			clk       : in std_logic;					  
			rst       : in std_logic;
		
	-- control signals from master controller.	
			mode      : in std_logic_vector(2 downto 0);
			op_1      : in std_logic_vector(3 downto 0);
			op_2      : in std_logic_vector(3 downto 0);
			op_r      : in std_logic_vector(3 downto 0);
		spec_command  : in std_logic_vector(2 downto 0);	-- certain modes has more options, and used to set special mast_ctrl functions.
		mat_order_in  : in std_logic_vector(5 downto 0);    -- to set the max value of registers that decide the order of the matrix.
	  dynamic_scale_in: in std_logic_vector(5 downto 0);
-- controls singals to mpma	
	m_muli_sel_reg    : out std_logic;                            -- mux at multiply inputs , active to select the register array.
    m_s1_adder_seli1  : out std_logic;     						  -- mux at the odd stage1 adder input1, 1 chooses the ram_data_in_1.
	m_s1_adder_seli2  : out std_logic_vector(1 downto 0);		  -- mux at the odd stage1 adder input2.
	m_data_out_sel    : out std_logic_vector(1 downto 0);         -- mux at the output stage.
                        
	s1_sub_e          : out std_logic;							  -- for add/ subtract operation.
    s1_acc_enable     : out std_logic;							  -- enable the accumulators at stage 1.
	s2_acc_enable     : out std_logic;							  -- enable the stage 2 accumulators
	flush             : out std_logic;                            -- to flush out the accumulators
	enc_dynamic_scale : out std_logic_vector(1 downto 0);         -- for dynamic scaling at the output. generated by master controller.

-- used for loading data in	
	i_data_vld        : in  std_logic;
    data_out_vld      : out std_logic;
	
-- control signals to address decoder.	
	ram_sel_out       : out  std_logic_vector(3 downto 0);
    write_en          : out  std_logic;
	row_cnt_out       : out  std_logic_vector(5 downto 0);
    row_set_out       : out  std_logic_vector(3 downto 0);
	mat_index_out     : out  std_logic_vector(3 downto 0);
-- control signals for register array.	
     row_i    		  : out  std_logic_vector(5 downto 0);		-- used to write to register array.
	 reg_rwn          : out  std_logic; 					    -- to read or write to register array.
   reg_row_set        : out  std_logic_vector(3 downto 0);      -- should be connected row_offset.
  
--
   data_in_sel        : out std_logic_vector(1 downto 0);
-- control signals for divider.
   div_row_mode       : out std_logic_vector(1 downto 0);
   div_address        : out std_logic_vector(7 downto 0) 
  
);
end entity;


architecture beh of mat_ctrl_v1 is

type system_state is (st_idle,							-- idle state.
														--used for loading matrix to RAM.
					  st_load_mat,
					  
					  st_load_mat_out,					-- used for loading matrix from RAM.
					  st_load_mat_out_wt,
														-- used for mat multiply.
					  st_load_row,						-- used to load 4 rows to register array.
					  st_load_row_wt,
					  st_read_ram,st_read_ram_wt,		-- used to read ram data.
					  st_write_ram,						    -- starts executing the current instruction.
					  st_s1_acc_update,					--used for mat_addi
							
														-- used for mat copy.
					  st_mc_read,						-- used for matrix  read.
                      st_mc_write,					    -- used for matrix write.
														-- used for matrix diag_add.
					  st_diag_add_read,
					  st_diag_add_write,
												
														--used for diagonal multiply operation
					 st_diag_mul_read,
                     st_diag_mul_write,					 
					 st_done);							-- reached the end of executing current instruction.

signal cs, ns   : system_state ;                		-- used for the state machine, next state and current state.

--- to make it work for all orders from 4 to 64.
signal rs_row_cnt_max,rs_row_cnt,
	   row_cnt_max,row_cnt, 
	   rs_row_cnt_incr,row_cnt_incr,
	   cs_reg_cnt,cs_reg_cnt_incr
						   : unsigned(5 downto 0);
signal row_set,row_set_max,
	   col_set,col_set_max,col_set_ff,
	   row_set_incr,col_set_incr,
	   reg_load_cnt,reg_load_cnt_max,
	   reg_load_cnt_incr,rs_row_set,
	   rs_row_set_incr
	                       : unsigned(3 downto 0);
						   
signal ram_sel,ram_sel_incr: unsigned(1 downto 0); --2 bits
signal ram_sel_all         : std_logic_vector(1 downto 0);
signal ram_sel_stored,
       ram_sel_stored_incr,
       rs_ram_sel,rs_ram_sel_incr
                    	   : unsigned(1 downto 0); -- used in matrix to matrix multiply to store the remsel value when leaving the load row state.

-- fix						   
--signal row_set_ff :  unsigned(3 downto 0);
						   
begin



--row_mode 01 for fetching same data over four outputs X*Z-1
--row_mode 10 for fetching different data from different location Z-1 *X
-- 
-- 
-- driving the divider addresses.
div_row_mode <="01" when spec_command ="000" else "10";
div_address  <= "00"&std_logic_vector(row_cnt) when spec_command ="000" 
                   else "00"&std_logic_vector(row_cnt(5 downto 2))&"00"; 


-- used for data mux at topdesign

 data_in_sel <= "00" when cs = st_load_mat else 
                "01" when cs = st_mc_read or cs = st_mc_write else
				"11"; -- for other operations.

--- used for the register array.

process(cs,row_cnt) 
begin
	if(cs =st_load_row or cs = st_load_row_wt) then
	   row_i <= std_logic_vector(row_cnt);
	 else
	   row_i <= (others =>'0');
	end if; 
	   
end process;

-- used 

process(cs)
begin
  if(cs = st_load_row or cs = st_load_row_wt) then
		reg_rwn <='0'; -- for writing.
  else
		reg_rwn <='1'; -- for reading.
  end if;

end process;


process(cs,col_set)
begin
 if(cs = st_read_ram or cs = st_read_ram_wt or cs = st_s1_acc_update
	or cs = st_write_ram) then
  reg_row_set <= std_logic_vector(col_set);
  else
   reg_row_set <=(others =>'0');
  end if;

end process;

-- used to select the mpma output mux.
process (cs) 
begin
	if(cs =st_diag_add_read or cs =st_diag_add_write) then
	 m_data_out_sel <="01";
	elsif(cs =st_diag_mul_read or cs= st_diag_mul_write) then
	 m_data_out_sel <= "10";
	else -- for matrix multiply operation.
	 m_data_out_sel <="00";
	end if; 
end process;

process(cs)
begin
    if(cs = st_diag_mul_read or cs =st_diag_mul_write) then
     m_muli_sel_reg <= '0' ;
    else -- to select data from register array.
     m_muli_sel_reg <='1';
    end if;
end process;

process(cs)
begin
	if(cs =st_diag_add_read or cs =st_diag_add_write) then
		m_s1_adder_seli1 <='0';
	else	-- matrix multiply.
		m_s1_adder_seli1 <='1';
	end if;
end process;

process(cs)
begin
	if(cs =st_diag_add_read or cs =st_diag_add_write) then
		m_s1_adder_seli2 <="01";
	else -- matrix multiply.
		m_s1_adder_seli2 <="00";	
	end if;
end process;


process(cs)
begin
	if(cs= st_done or cs = st_write_ram or cs = st_idle)then -- just to make sure the accumulators are clean.
	   flush <='1';
	else
	   flush <='0';
	end if;  
end process; 

  
process(cs, spec_command) begin
	if((cs = st_diag_add_read or cs= st_diag_add_write)and spec_command="001") then     
		s1_sub_e <='1';		-- do subtract.
	else
		s1_sub_e <='0';		-- do addition.
	end if; 
end process;

process(cs) begin
	if(cs= st_s1_acc_update) then
	  s1_acc_enable <='1';
	else
	  s1_acc_enable <='0';  
	end if;  
end process;

          
--dynamic_scale   , driven by master controller based on instruction. no encoding needed  for now.
-- dynamic scale encoder




-- only need to generate for the  dynamic scale needed. but for the general case, I am splitting the dynamic scale into four sections to 
-- reduce the size of MUX at the ouput stage od PMPA.
process(dynamic_scale_in)
 begin
	   if(dynamic_scale_in < "010000") then -- less than 16
	  enc_dynamic_scale <= "00";
	elsif(dynamic_scale_in < "100000") then	-- less than 32
	  enc_dynamic_scale <= "01";
	elsif(dynamic_scale_in < "110000") then -- less than 48
	  enc_dynamic_scale <= "10";
	else                                    -- less than 64.
	  enc_dynamic_scale <= "11";
	end if;
end process;

   
--s2_acc_enable   to be used only for mat to mat addition and mat to mat dot product. not  implemented for the Matrix inverse.
s2_acc_enable <='0';


--- used to drive the address decoder.

row_cnt_out_gen: process(row_cnt,rs_row_cnt,cs)
begin

	if( cs = st_write_ram or cs = st_read_ram or cs = st_read_ram_wt or cs = st_s1_acc_update) then
		row_cnt_out <= std_logic_vector(rs_row_cnt);
	else
        row_cnt_out <= std_logic_vector(row_cnt);
	end if;


end process;





-- selecting the row set based on the operation.
row_set_out_gen : process(row_set,col_set,cs,rs_row_set)
begin
  if(cs =st_read_ram or cs = st_read_ram_wt or cs= st_s1_acc_update) then		
       row_set_out <= std_logic_vector(col_set);
  elsif(cs = st_write_ram or cs = st_load_row or cs= st_load_row_wt) then
       row_set_out <= std_logic_vector(rs_row_set);  
  else
	   row_set_out <= std_logic_vector(row_set);
  end if;

end process; 

-- generate the right index for the matrix.
mat_index_out_gen: process(op_1,op_2,op_r,cs)
begin

	if(  cs = st_mc_read or cs = st_diag_mul_read or 
		 cs = st_load_row or cs = st_load_row_wt)then
		mat_index_out <= op_1;
	elsif(cs = st_read_ram or cs= st_read_ram_wt or cs =st_s1_acc_update) then
		mat_index_out <= op_2;
	else-- rest of the states uses op_r.
		mat_index_out <= op_r;
	end if;


end process;







--- used when all of the ram are read or write.
ram_sel_all <= "01" when cs = st_diag_mul_read or cs = st_diag_mul_write or
						 cs = st_read_ram or cs = st_read_ram_wt or 
						 cs = st_s1_acc_update or cs = st_mc_read or cs= st_mc_write or
                         cs = st_read_ram or cs= st_read_ram_wt						 else -- to select all ram.
			   "10" when cs = st_idle												 else -- to deselect all ram.
			   "00" ;
			   
			   
-- ram_sel out generator.			   
process (ram_sel_all, ram_sel,cs,row_cnt,ram_sel_stored,rs_ram_sel )
begin

if(cs =st_diag_add_read or cs= st_diag_add_write )  then		        -- for diagonal addition operation.
	 ram_sel_out <= ram_sel_all& std_logic_vector(row_cnt(1 downto 0)); -- used for mat to diag matrix addition.

elsif(cs = st_load_row or cs = st_load_row_wt) then 					-- used for loading the register to the ROW.
     ram_sel_out <= ram_sel_all & std_logic_vector(ram_sel_stored);
elsif(cs = st_write_ram) then
     ram_sel_out <=	ram_sel_all & std_logic_vector(rs_ram_sel);
else
	 ram_sel_out <= ram_sel_all & std_logic_vector(ram_sel); 			-- generate the ram_sel signal for address decoder.
end if;
end process;

-- write enable is set to 1 when cs= st_mc_write or cs = st_load_mat
write_en    <= '1' when cs= st_load_mat or cs = st_diag_mul_write
						or cs = st_mc_write or cs = st_load_mat     -- enable write to RAM.
						or cs = st_diag_add_write or cs = st_write_ram
		  else '0';
		  
-- data out valid when cs is st_load_mat_out_wt
data_out_vld  <= '1' when cs = st_load_mat_out_wt else '0';

  

-- for now only square matrices are considered.
-- controls how long the states are performed.
process (mat_order_in)
begin
	rs_row_cnt_max   <= unsigned(mat_order_in)-1;
	row_cnt_max      <= unsigned(mat_order_in)-1;
	col_set_max      <= unsigned(mat_order_in(5 downto 2))-1;
	row_set_max      <= unsigned(mat_order_in(5 downto 2))-1;
	reg_load_cnt_max <= unsigned(mat_order_in(5 downto 2))-1;
end process;


-- ram_sel increment to switch to the next ram .

ram_sel_incr_gen: process(cs,row_cnt,row_cnt_max,
						  ram_sel
						 )
begin
	if((cs= st_load_mat and row_cnt = row_cnt_max)         or
	    (cs= st_load_mat_out_wt and row_cnt = row_cnt_max) or 
		(cs = st_write_ram)
	  ) then
	      
					ram_sel_incr <= ram_sel +1;
		  
	--elsif(cs =st_diag_add_read or cs= st_diag_add_write )  then		-- for diagonal addition operation.
	 -- ram_sel_incr <= row_cnt(1 downto 0); doesn't work this way, have to mux the ram_sel out 
	else
	  ram_sel_incr <= ram_sel;
	end if;  
end process; 


--store ram_Sel value. used for loading row data into register.

ram_sel_stored_incr_gen: process(cs,ram_sel_stored,row_cnt_max,row_cnt)

begin
if(cs = st_load_row_wt and row_cnt = row_cnt_max) then
	 ram_sel_stored_incr <= ram_sel_stored+1;		-- store the ram_sel here.
else
     ram_sel_stored_incr <= ram_sel_stored;
end if;

end process;


--- generate to navigate the elements of the row..
row_cnt_incr_gen: process(cs,row_cnt,i_data_vld,row_cnt_max)
begin
	 if((cs= st_load_mat and i_data_vld='1') or   -- for loading matrix in.
			cs = st_load_mat_out_wt or			  -- for loading matrix out.
			cs = st_mc_write	or				  -- for matrix copy.
			cs = st_load_row_wt or 				  -- for matrix multiply
			cs = st_diag_mul_write or			  -- for matrix diagonal multiply
			cs = st_diag_add_write 				  -- for matrix diagonal addition.
			
			
		) then				  
		   if(row_cnt=row_cnt_max) then	
				row_cnt_incr <= (others=>'0');
		   else
				row_cnt_incr <= row_cnt+1;
		   end if;		   
	 
	 elsif(cs = st_done and row_cnt= row_cnt_max) then
	       row_cnt_incr <= (others=>'0');
	 else
	 
		row_cnt_incr <= row_cnt;
	 end if;

end process;

-- used to goto next set of rows in the RAM.
row_set_incr_gen: process(cs,row_set,row_cnt,row_cnt_max,row_set_max,
						  ram_sel)
begin
	 if((cs= st_load_row_wt and ram_sel="11") or
	    (cs= st_diag_mul_write and row_cnt= row_cnt_max) or
		(cs= st_mc_write and row_cnt = row_cnt_max) or
		((cs = st_load_mat or cs = st_load_mat_out_wt) and row_cnt = row_cnt_max and ram_sel="11") or
		(cs = st_diag_add_write and row_cnt(1 downto 0)="11")
		)then
		if(row_set=row_set_max) then		
			row_set_incr<="0000";		-- clears to one if it reaches the max point.
		else
			row_set_incr <= row_set+1;			-- increments rowset.
		end if;
	     
		 
		 
	 else
		row_set_incr <= row_set;
	 end if;

end process;



-- used during the st_ram_write stage. for writing results during the RAM write state.
rs_row_cnt_incr_gen: process(cs,rs_row_cnt, row_cnt_max)
begin
	if(cs=st_write_ram) then -- get the next row into ram.
		if(rs_row_cnt = row_cnt_max) then
			rs_row_cnt_incr <= (others=>'0'); 
		else
			rs_row_cnt_incr <= rs_row_cnt +1;
		end if;
		
	else
		rs_row_cnt_incr <= rs_row_cnt;
	end if;
end process;

rs_row_set_incr_gen : process(rs_row_set,rs_ram_sel,row_set_max,
							  cs,rs_row_cnt,row_cnt_max	)
begin
	if(rs_ram_sel="11" and rs_row_cnt= row_cnt_max and cs = st_write_ram) then
		if(rs_row_set = row_set_max) then
		    rs_row_set_incr <= (others=>'0');
		else
		    rs_row_set_incr <= rs_row_set +1;
		end if;
	else
			rs_row_set_incr <= rs_row_set; 
	end if;

end process;




rs_ram_sel_gen : process(rs_row_cnt,row_cnt_max,cs,rs_ram_sel)
begin
	if(rs_row_cnt=row_cnt_max and cs = st_write_ram) then
	 rs_ram_sel_incr <= rs_ram_sel+1;
	else
	 rs_ram_sel_incr <= rs_ram_sel;
	end if;
end process;




---

cs_reg_cnt_gen: process(cs, cs_reg_cnt,row_cnt_max,ns)
begin
 if(ns= st_read_ram and cs = st_load_row_wt) then	-- during the transaction to row to mat multiply stage.
    if(cs_reg_cnt= row_cnt_max) then
	    cs_reg_cnt_incr <= (others =>'0');
	else
		cs_reg_cnt_incr <= cs_reg_cnt+1;
	end if;
 elsif(cs = st_done) then
    cs_reg_cnt_incr <= (others =>'0');
 else
    cs_reg_cnt_incr <= cs_reg_cnt;
 end if;
end process;


col_set_incr_gen: process(cs,col_set,col_set_max) 
begin
	if(cs= st_read_ram_wt) then
		 if(col_set=col_set_max) then		
				col_set_incr<="0000";		-- clears to one if it reaches the max point.
			else
				col_set_incr <= col_set+1;			-- increments colset.
			end if;
		 else
			col_set_incr <= col_set;
    end if;

end process;



done <= '1' when cs= st_done else '0';


--- the registers used to drive the mat controller. 

statemachine_seq: process(clk,rst)
begin
if(rst='1') then
					cs  <=  st_idle;
			 rs_row_cnt <= (others=>'0');
				row_cnt <= (others=>'0');
				col_set <= (others=>'0');
				row_set <= (others=>'0'); 
				ram_sel <= (others=>'0');
		 ram_sel_stored <= (others=>'0');
             rs_row_set <= (others=>'0');
			 rs_ram_sel <= (others=>'0');
			 cs_reg_cnt <= (others=>'0');
			 col_set_ff <= (others=>'0');
		--	 row_set_ff <= (others=>'0');
elsif(rising_edge(clk)) then
					cs  <= ns;
		     rs_row_cnt <= rs_row_cnt_incr;
			 rs_ram_sel <= rs_ram_sel_incr;
			 rs_row_set <= rs_row_set_incr;
				row_cnt <= row_cnt_incr;
				col_set <= col_set_incr;
				row_set <= row_set_incr;
				ram_sel <= ram_sel_incr;
		 ram_sel_stored <= ram_sel_stored_incr;
		     cs_reg_cnt <= cs_reg_cnt_incr;
			 col_set_ff <= col_set;
			-- row_set_ff <= row_set;
end if;
end process;



-- state machine for all the operations supported for now./

statemachine_comb: process(cs, start,
							ram_sel, row_cnt,row_cnt_max,
							rs_row_cnt,rs_row_cnt_max,col_set,
							col_set_max,mode,col_set_ff,
							row_set,row_set_max,cs_reg_cnt,rs_ram_sel,
							rs_row_set)
begin
	case cs is
	 when st_idle =>
		 if(start='1') then
		    case mode is	 -- branches to different state machines.
			 when "000" =>   -- matrix load to RAM
				ns <= st_load_mat;
			 when "001" =>   -- matrix to matrix multipication.
				ns <= st_load_row;
			 when "100" =>   --matrix copy.	
			    ns <= st_mc_read;
			 when "010" =>	 -- diag mulitplication. 
                ns <= st_diag_mul_read;
             when "011" =>   -- diag_addition.
                ns <= st_diag_add_read;			 
			 when "111" =>
				ns <= st_load_mat_out;
			 when others =>
				ns <= st_idle; 	 
		    end case;		
		 else
		  ns <= st_idle;
		 end if;
		 
-- for matrix load operation in .		 
     when st_load_mat=>
        if(ram_sel= "11" and row_cnt= row_cnt_max and row_set = row_set_max) then
		  ns <= st_done; --- reached the end of writing.
		else
		  ns <= st_load_mat;
		end if;
-- for matrix load out operation.
     when st_load_mat_out =>
	    ns <= st_load_mat_out_wt;
	 when st_load_mat_out_wt =>
	    if(ram_sel= "11" and row_cnt= row_cnt_max and row_set = row_set_max) then
		  ns <= st_done; --- reached the end of reading.
		else
		  ns <= st_load_mat_out;
		end if;
-- for matrix copy		
     when st_mc_read  =>
		ns <= st_mc_write;
	 when st_mc_write =>
   	    if(row_set=row_set_max and row_cnt= row_cnt_max) then
		  ns <= st_done; --- reached the end of writing.
		else
		  ns <= st_mc_read;
		end if;
--	for diag mulitplication
     when st_diag_mul_read =>
	      ns <= st_diag_mul_write;
	 when st_diag_mul_write =>
	    if(row_set= row_set_max and row_cnt= row_cnt_max) then
		  ns <= st_done; --- reached the end of writing.
		else
		  ns <= st_diag_mul_read;
		end if;
--  for diag_ addition operation		
	  when st_diag_add_read  =>
		  ns <= st_diag_add_write;
	  when st_diag_add_write =>
		  if(row_cnt= row_cnt_max) then
		   ns <= st_done;
		  else
		   ns <= st_diag_add_read;
		  end if;
-- for matrix multiply operation	 
	 -- loading register arrays with 4 rows from RAM.
	 when st_load_row=>
	   ns <= st_load_row_wt;
	 when st_load_row_wt =>	   
	  if(row_cnt= row_cnt_max) then	
	   ns <= st_read_ram;		--update row_set by 1 
	  else
	   ns <= st_load_row;
	  end if;
	  -- starting matrix multiply with the current set of 4 rows. 
	 when st_read_ram =>
	  ns<= st_read_ram_wt;
	 when st_read_ram_wt=>
      
	    if(col_set=(col_set_max)) then -- the last step should be st_write_ram
		   ns <= st_write_ram; -- at the end of last set of matrix.
		  else
		   ns <= st_s1_acc_update;
		  end if;
	 when st_s1_acc_update=> 
	     ns <= st_read_ram_wt;
			
     when st_write_ram =>
	   if(ram_sel= "11" and col_set_ff = col_set_max and 
		    rs_row_cnt=rs_row_cnt_max) then -- found result for one row of resultant matrix.
														-- increment row_cnt.
														-- load the ramsel_stored back to ram_sel.
														-- increment col_set.
			--if(rs_ram_sel="11" and rs_row_set= row_set_max) then -- found results for the last row. check rs_row_set and rs_ram_sel
			if(cs_reg_cnt="000000" and rs_ram_sel="11" and rs_row_set=row_set_max) then
			  ns <= st_done;
			else
			  ns <= st_load_row;
			end if;
	   else
		 ns <= st_read_ram;
	   end if;
     when st_done =>
      ns <= st_idle;	 
	  -- generate ok handshake to end the current executing.
	 when  others=>
	  ns <= st_idle;
	end case;

end process;


end beh;